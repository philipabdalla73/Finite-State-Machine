LIBRARY ieee ;
USE ieee.std_logic_1164.all ;
ENTITY SSEG IS
PORT ( bcd : IN STD_LOGIC_VECTOR(3 DOWNTO 0) ;
Sign : IN STD_LOGIC;
leds : OUT STD_LOGIC_VECTOR(1 TO 7);
ledss : OUT STD_LOGIC_VECTOR(1 TO 7));
END SSEG;

ARCHITECTURE Behavior OF SSEG IS
BEGIN
PROCESS ( bcd )
BEGIN
CASE bcd IS          -- abcdefg
WHEN "0000" => leds <= "0000001";--0
WHEN "0001" => leds <= "1111001";--1
WHEN "0010" => leds <= "0010010";--2
WHEN "0011" => leds <= "0000110";--3
WHEN "0100" => leds <= "1001100";--4
WHEN "0101" => leds <= "0100100";--5
WHEN "0110" => leds <= "0100000";--6
WHEN "0111" => leds <= "0001111";--7
WHEN "1000" => leds <= "0000000";--8
WHEN "1001" => leds <= "0001100";--9


WHEN "1010" => leds <= "0001000";--10
WHEN "1011" => leds <= "1100000";--11
WHEN "1100" => leds <= "0110001";--12
WHEN "1101" => leds <= "1000010";--13
WHEN "1110" => leds <= "0110000";--14
WHEN "1111" => leds <= "0111000";--15
WHEN OTHERS => leds <= "-------" ;
END CASE ;
CASE Sign IS       -- abcdefg
WHEN '1' => ledss <= "1111110";
WHEN '0' => ledss <= "1111111";
WHEN OTHERS => leds <= "-------" ;
END CASE ;
END PROCESS ;
END Behavior ;